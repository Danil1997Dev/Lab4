 

module sdmodb 
(
    input clk,clr_n,
	 input signed [7:0] val,// входные данные модулятора; 
	 output daco //однобитная выходная последовательность.
); 
  
  reg signed [7:0] daco_reg = 0;
  reg signed [7:0] val_delay = 0;
  reg signed [7:0] val_def = 0;
  reg signed [7:0] val_delay_compar = 0;

  always @(posedge clk or negedge clr_n)
    begin
      if (!clr_n)
        begin
			  daco_reg  = 1'b0;
			  val_delay = 1'b0;
        end
      else
        begin
			val_def = val - daco_reg;
			val_delay <= val_def + val_delay;
			val_delay_compar <= val_delay;
			if (val_delay >= val_delay_compar) begin
			  daco_reg =  127;  end
			else begin
			  daco_reg = -127;  end
        end
    end 
	
  assign daco = daco_reg[7];
  
endmodule

