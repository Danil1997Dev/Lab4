
module niosII (
	clk_clk,
	reset_reset_n,
	generator_export_fout);	

	input		clk_clk;
	input		reset_reset_n;
	output		generator_export_fout;
endmodule
